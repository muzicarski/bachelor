`ifndef __BRAM_UVM_PKG_SV__
`define __BRAM_UVM_PKG_SV__

package bram_uvm_pkg;

   import uvm_pkg::*;
`include "uvm_macros.svh"

`include "bram_monitor.sv"
   
   
endpackage // bram_uvm_pkg

`endif
   
